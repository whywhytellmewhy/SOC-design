// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none

`timescale 1 ns / 1 ps

module counter_la_fir_tb;
	reg clock;
        reg RSTB;
	reg CSB;

	reg power1, power2;

	wire gpio;
	wire uart_tx;
	wire [37:0] mprj_io;
	wire [15:0] checkbits;

	assign checkbits  = mprj_io[31:16];
	assign uart_tx = mprj_io[6];

	always #12.5 clock <= (clock === 1'b0);

	initial begin
		clock = 0;
	end

	`ifdef ENABLE_SDF
		initial begin
			$sdf_annotate("../../../sdf/user_proj_example.sdf", uut.mprj) ;
			$sdf_annotate("../../../sdf/user_project_wrapper.sdf", uut.mprj.mprj) ;
			$sdf_annotate("../../../mgmt_core_wrapper/sdf/DFFRAM.sdf", uut.soc.DFFRAM_0) ;
			$sdf_annotate("../../../mgmt_core_wrapper/sdf/mgmt_core.sdf", uut.soc.core) ;
			$sdf_annotate("../../../caravel/sdf/housekeeping.sdf", uut.housekeeping) ;
			$sdf_annotate("../../../caravel/sdf/chip_io.sdf", uut.padframe) ;
			$sdf_annotate("../../../caravel/sdf/mprj_logic_high.sdf", uut.mgmt_buffers.mprj_logic_high_inst) ;
			$sdf_annotate("../../../caravel/sdf/mprj2_logic_high.sdf", uut.mgmt_buffers.mprj2_logic_high_inst) ;
			$sdf_annotate("../../../caravel/sdf/mgmt_protect_hv.sdf", uut.mgmt_buffers.powergood_check) ;
			$sdf_annotate("../../../caravel/sdf/mgmt_protect.sdf", uut.mgmt_buffers) ;
			$sdf_annotate("../../../caravel/sdf/caravel_clocking.sdf", uut.clocking) ;
			$sdf_annotate("../../../caravel/sdf/digital_pll.sdf", uut.pll) ;
			$sdf_annotate("../../../caravel/sdf/xres_buf.sdf", uut.rstb_level) ;
			$sdf_annotate("../../../caravel/sdf/user_id_programming.sdf", uut.user_id_value) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_bidir_1[0] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_bidir_1[1] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_bidir_2[0] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_bidir_2[1] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_bidir_2[2] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_1[0] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_1[1] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_1[2] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_1[3] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_1[4] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_1[5] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_1[6] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_1[7] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_1[8] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_1[9] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_1[10] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_1a[0] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_1a[1] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_1a[2] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_1a[3] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_1a[4] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_1a[5] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_2[0] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_2[1] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_2[2] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_2[3] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_2[4] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_2[5] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_2[6] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_2[7] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_2[8] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_2[9] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_2[10] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_2[11] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_2[12] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_2[13] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_2[14] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_control_block.sdf", uut.\gpio_control_in_2[15] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.\gpio_defaults_block_0[0] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.\gpio_defaults_block_0[1] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.\gpio_defaults_block_2[0] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.\gpio_defaults_block_2[1] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.\gpio_defaults_block_2[2] ) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_5) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_6) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_7) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_8) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_9) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_10) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_11) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_12) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_13) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_14) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_15) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_16) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_17) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_18) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_19) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_20) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_21) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_22) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_23) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_24) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_25) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_26) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_27) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_28) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_29) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_30) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_31) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_32) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_33) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_34) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_35) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_36) ;
			$sdf_annotate("../../../caravel/sdf/gpio_defaults_block.sdf", uut.gpio_defaults_block_37) ;
		end
	`endif 

	// assign mprj_io[3] = 1'b1;

	initial begin
		$dumpfile("counter_la_fir.vcd");
		$dumpvars(0, counter_la_fir_tb);

		// Repeat cycles of 1000 clock edges as needed to complete testbench
		repeat (2500) begin // modified (original:250)
			repeat (1000) @(posedge clock);
			// $display("+1000 cycles");
		end
		$display("%c[1;31m",27);
		`ifdef GL
			$display ("Monitor: Timeout, Test LA (GL) Failed");
		`else
			$display ("Monitor: Timeout, Test LA (RTL) Failed");
		`endif
		$display("%c[0m",27);
		$finish;
	end

	initial begin
		wait(checkbits == 16'hAB40);
		$display("LA Test 1 started");
		//wait(checkbits == 16'hAB41);

		//wait(checkbits == 16'd40);
		//$display("Call function matmul() in User Project BRAM (mprjram, 0x38000000) return value passed, 0x%x", checkbits);
		//wait(checkbits == 16'd893);
		//$display("Call function matmul() in User Project BRAM (mprjram, 0x38000000) return value passed, 0x%x", checkbits);
		//wait(checkbits == 16'd2541);
		//$display("Call function matmul() in User Project BRAM (mprjram, 0x38000000) return value passed, 0x%x", checkbits);
		//wait(checkbits == 16'd2669);
		//$display("Call function matmul() in User Project BRAM (mprjram, 0x38000000) return value passed, 0x%x", checkbits);		

		///////////////////////////////// Added /////////////////////////////////
		/*wait(checkbits == 16'd10614); //////////////////////<----------------------------------------------------- remember to uncomment this !!!!!
		$display("Call \"software\" function fir() in User Project BRAM (mprjram, 0x38000000) return value passed, 0x%x, which is %d in decimal", checkbits, checkbits);
		*/
		/////wait(checkbits == 16'd123);
		/////$display("Call function fir() in User Project BRAM (mprjram, 0x38000000) return value passed, 0x%x, which is %d in decimal", checkbits, checkbits);
		/////////////////////////////////////////////////////////////////////////
		
		wait(checkbits == 16'hAB51);
		$display("LA Test 2 passed");

		///////////////////////////////// Added /////////////////////////////////
		$display("---------------------------------------------");
        $display("-----------Congratulations! Pass-------------");
		/////////////////////////////////////////////////////////////////////////

		#10000;
		$finish;
	end

	// Added by us to assist notification when some error happens
	initial begin
		//wait(checkbits == 16'hFFFF);
		//$display("Error: Something wrong, so fir.c returned \"-1\" !!!");
		wait(checkbits == 16'hFFFE);
		$display("Error: Something wrong, so fir.c returned \"-2\" !!!");
		$display("--------Simulation Failed---------");
		#10000;
		$finish;
	end
	// Added by us to assist notification when some error happens
	initial begin
		wait(checkbits == 16'hFFFD);
		$display("Error: Something wrong, so fir.c returned \"-3\" !!!");
		$display("--------Simulation Failed---------");
		#10000;
		$finish;
	end

	// Added by us to build a latency_timer
	integer latency_timer;
    initial begin
        latency_timer = 0;
        #5;
        forever begin
            #10 latency_timer = latency_timer+1;
        end
    end

	// Added by us to count latency_timer
	integer FIR_latency_firmware;
	integer FIR_latency_round1;
	integer FIR_latency_round2;
	integer FIR_latency_round3;
	integer golden_final_Y;
	initial begin
		golden_final_Y=10614;
		///////////////////////////////////// For firmware /////////////////////////////////////
		$display("\n++++++++++ Step 1: Use firmware (lab4-1) ++++++++++");
		wait(checkbits[7:0] == 8'hA5);
		latency_timer=0;
		$display("(Firmware) Detect start mark (8'hA5) on mprj[23:16], start latency timer.");
		wait(checkbits[7:0] == 8'h5A);
		FIR_latency_firmware=latency_timer;
		$display("(Firmware) Detect end mark (8'h5A) on mprj[23:16], record latency timer.");
		if (checkbits[15:8] == golden_final_Y[7:0]) begin
			$display("(Firmware) Success: Final Y[7:0] output to mprj[31:24] is 0x%x, the same as the golden value.", checkbits[15:8]);
		end
		else begin
			$display("(Firmware) Error: Final Y[7:0] output to mprj[31:24] is 0x%x, which is NOT the same as the golden value.", checkbits[15:8]);
			$display("--------Simulation Failed---------");
			$finish;
		end
        $display("Info: FIR \"firmware\" latency = %d clock cycles", FIR_latency_firmware);

		$display("\n++++++++++ Step 2: Use hardware (FIR engine)(lab3) ++++++++++");
		///////////////////////////////////// For round 1 /////////////////////////////////////
		wait(checkbits[7:0] == 8'hA5);
		latency_timer=0;
		$display("(Round 1) Detect start mark (8'hA5) on mprj[23:16], start latency timer.");
		wait(checkbits[7:0] == 8'h5A);
		FIR_latency_round1=latency_timer;
		$display("(Round 1) Detect end mark (8'h5A) on mprj[23:16], record latency timer.");
		///// 5. compare Yn with golden data (lab3 workbook p.19)
        ///// 3. Checking phase: (2)Compare Yn buffer with golden data (lab3 workbook p.20)
		/////if (checkbits[15:8] == 8'd10614) begin
		if (checkbits[15:8] == golden_final_Y[7:0]) begin
			$display("(Round 1) Success: Final Y[7:0] output to mprj[31:24] is 0x%x, the same as the golden value.", checkbits[15:8]);
		end
		else begin
			$display("(Round 1) Error: Final Y[7:0] output to mprj[31:24] is 0x%x, which is NOT the same as the golden value.", checkbits[15:8]);
			$display("--------Simulation Failed---------");
			$finish;
		end
		///// 3. Checking phase: (1)Report latency (lab3 workbook p.20)
        $display("Info: FIR engine (hardware) latency in round 1 = %d clock cycles", FIR_latency_round1);

		///////////////////////////////////// For round 2 /////////////////////////////////////
		wait(checkbits[7:0] == 8'hA5);
		latency_timer=0;
		$display("(Round 2) Detect start mark (8'hA5) on mprj[23:16], start latency timer.");
		wait(checkbits[7:0] == 8'h5A);
		FIR_latency_round2=latency_timer;
		$display("(Round 2) Detect end mark (8'h5A) on mprj[23:16], record latency timer.");
		///// 5. compare Yn with golden data (lab3 workbook p.19)
        ///// 3. Checking phase: (2)Compare Yn buffer with golden data (lab3 workbook p.20)
		/////if (checkbits[15:8] == 8'd10614) begin
		if (checkbits[15:8] == golden_final_Y[7:0]) begin
			$display("(Round 2) Success: Final Y[7:0] output to mprj[31:24] is 0x%x, the same as the golden value.", checkbits[15:8]);
		end
		else begin
			$display("(Round 2) Error: Final Y[7:0] output to mprj[31:24] is 0x%x, which is NOT the same as the golden value.", checkbits[15:8]);
			$display("--------Simulation Failed---------");
			$finish;
		end
		///// 3. Checking phase: (1)Report latency (lab3 workbook p.20)
        $display("Info: FIR engine (hardware) latency in round 2 = %d clock cycles", FIR_latency_round2);

		///////////////////////////////////// For round 3 /////////////////////////////////////
		wait(checkbits[7:0] == 8'hA5);
		latency_timer=0;
		$display("(Round 3) Detect start mark (8'hA5) on mprj[23:16], start latency timer.");
		wait(checkbits[7:0] == 8'h5A);
		FIR_latency_round3=latency_timer;
		$display("(Round 3) Detect end mark (8'h5A) on mprj[23:16], record latency timer.");
		///// 5. compare Yn with golden data (lab3 workbook p.19)
        ///// 3. Checking phase: (2)Compare Yn buffer with golden data (lab3 workbook p.20)
		/////if (checkbits[15:8] == 8'd10614) begin
		if (checkbits[15:8] == golden_final_Y[7:0]) begin
			$display("(Round 3) Success: Final Y[7:0] output to mprj[31:24] is 0x%x, the same as the golden value.", checkbits[15:8]);
		end
		else begin
			$display("(Round 3) Error: Final Y[7:0] output to mprj[31:24] is 0x%x, which is NOT the same as the golden value.", checkbits[15:8]);
			$display("--------Simulation Failed---------");
			$finish;
		end
		///// 3. Checking phase: (1)Report latency (lab3 workbook p.20)
        $display("Info: FIR engine (hardware) latency in round 3 = %d clock cycles", FIR_latency_round3);

		$display("Info: Total FIR engine (hardware) latency = %d clock cycles", FIR_latency_round1+FIR_latency_round2+FIR_latency_round3);
	end

	initial begin
		RSTB <= 1'b0;
		CSB  <= 1'b1;		// Force CSB high
		#2000;
		RSTB <= 1'b1;	    	// Release reset
		#170000;
		CSB = 1'b0;		// CSB can be released
	end

	initial begin		// Power-up sequence
		power1 <= 1'b0;
		power2 <= 1'b0;
		#200;
		power1 <= 1'b1;
		#200;
		power2 <= 1'b1;
	end

	wire flash_csb;
	wire flash_clk;
	wire flash_io0;
	wire flash_io1;

	wire VDD1V8;
	wire VDD3V3;
	wire VSS;
    
	assign VDD3V3 = power1;
	assign VDD1V8 = power2;
	assign VSS = 1'b0;

	assign mprj_io[3] = 1;  // Force CSB high.
	assign mprj_io[0] = 0;  // Disable debug mode

	caravel uut (
/*
		.vddio	  (VDD3V3),
		.vddio_2  (VDD3V3),
		.vssio	  (VSS),
		.vssio_2  (VSS),
		.vdda	  (VDD3V3),
		.vssa	  (VSS),
		.vccd	  (VDD1V8),
		.vssd	  (VSS),
		.vdda1    (VDD3V3),
		.vdda1_2  (VDD3V3),
		.vdda2    (VDD3V3),
		.vssa1	  (VSS),
		.vssa1_2  (VSS),
		.vssa2	  (VSS),
		.vccd1	  (VDD1V8),
		.vccd2	  (VDD1V8),
		.vssd1	  (VSS),
		.vssd2	  (VSS),
*/
		.clock    (clock),
		.gpio     (gpio),
		.mprj_io  (mprj_io),
		.flash_csb(flash_csb),
		.flash_clk(flash_clk),
		.flash_io0(flash_io0),
		.flash_io1(flash_io1),
		.resetb	  (RSTB)
	);

	spiflash #(
		.FILENAME("counter_la_fir.hex")
	) spiflash (
		.csb(flash_csb),
		.clk(flash_clk),
		.io0(flash_io0),
		.io1(flash_io1),
		.io2(),			// not used
		.io3()			// not used
	);

	// Testbench UART
	tbuart tbuart (
		.ser_rx(uart_tx)
	);

endmodule
`default_nettype wire
